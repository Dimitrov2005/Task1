module phy(
	   input
	   in1,
	   in2,
	   in3,
	   output reg
	   out1,
	   out2,
	   out3
	   );
   
   assign out1='bx;
   assign out2='bx;
   assign out3='bx;
   
endmodule // phy
