interface iface(input logic TCLK,TRESETN);
   logic TMS, 
	 WSI,
	 WSO;
endinterface